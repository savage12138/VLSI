* SPICE NETLIST
***************************************

.SUBCKT TAPCELL
** N=4 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_1
** N=6 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT M1_N_CDNS_586572660572
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT M1_POLY_CDNS_586572660570
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT M2_M1_via
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT M1_P_CDNS_586572660571
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_2
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT FullAdderMirror CIN VDD A B COUT GND SUM
** N=23 EP=7 IP=57 FDC=28
M0 GND A 10 GND NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.07e-14 PD=6.4e-07 PS=5.9e-07 $X=390 $Y=355 $D=1
M1 21 A GND GND NMOS_VTL L=5e-08 W=1.8e-07 AD=2.565e-14 AS=2.52e-14 PD=6.45e-07 PS=6.4e-07 $X=770 $Y=355 $D=1
M2 11 B 21 GND NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.565e-14 PD=6.4e-07 PS=6.45e-07 $X=1155 $Y=355 $D=1
M3 10 CIN 11 GND NMOS_VTL L=5e-08 W=1.8e-07 AD=2.565e-14 AS=2.52e-14 PD=6.45e-07 PS=6.4e-07 $X=1535 $Y=355 $D=1
M4 GND B 10 GND NMOS_VTL L=5e-08 W=1.8e-07 AD=3.15e-14 AS=2.565e-14 PD=8.2e-07 PS=6.45e-07 $X=1920 $Y=355 $D=1
M5 22 B GND GND NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=3.15e-14 PD=8.2e-07 PS=8.2e-07 $X=2300 $Y=175 $D=1
M6 23 A 22 GND NMOS_VTL L=5e-08 W=2.7e-07 AD=3.8475e-14 AS=3.78e-14 PD=8.25e-07 PS=8.2e-07 $X=2680 $Y=175 $D=1
M7 13 CIN 23 GND NMOS_VTL L=5e-08 W=2.7e-07 AD=3.15e-14 AS=3.8475e-14 PD=8.2e-07 PS=8.25e-07 $X=3065 $Y=175 $D=1
M8 15 11 13 GND NMOS_VTL L=5e-08 W=1.8e-07 AD=2.565e-14 AS=3.15e-14 PD=6.45e-07 PS=8.2e-07 $X=3445 $Y=355 $D=1
M9 GND CIN 15 GND NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.565e-14 PD=6.4e-07 PS=6.45e-07 $X=3830 $Y=355 $D=1
M10 15 A GND GND NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=4210 $Y=355 $D=1
M11 GND B 15 GND NMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.52e-14 PD=5.9e-07 PS=6.4e-07 $X=4590 $Y=355 $D=1
M12 COUT 11 GND GND NMOS_VTL L=5e-08 W=9e-08 AD=1.035e-14 AS=1.035e-14 PD=4.1e-07 PS=4.1e-07 $X=5450 $Y=535 $D=1
M13 SUM 13 GND GND NMOS_VTL L=5e-08 W=9e-08 AD=1.035e-14 AS=1.035e-14 PD=4.1e-07 PS=4.1e-07 $X=6310 $Y=535 $D=1
M14 VDD A 12 VDD PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=4.14e-14 PD=1e-06 PS=9.5e-07 $X=390 $Y=1960 $D=0
M15 18 A VDD VDD PMOS_VTL L=5e-08 W=3.6e-07 AD=5.13e-14 AS=5.04e-14 PD=1.005e-06 PS=1e-06 $X=770 $Y=1960 $D=0
M16 11 B 18 VDD PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=5.13e-14 PD=1e-06 PS=1.005e-06 $X=1155 $Y=1960 $D=0
M17 12 CIN 11 VDD PMOS_VTL L=5e-08 W=3.6e-07 AD=5.13e-14 AS=5.04e-14 PD=1.005e-06 PS=1e-06 $X=1535 $Y=1960 $D=0
M18 VDD B 12 VDD PMOS_VTL L=5e-08 W=3.6e-07 AD=6.3e-14 AS=5.13e-14 PD=1.36e-06 PS=1.005e-06 $X=1920 $Y=1960 $D=0
M19 19 B VDD VDD PMOS_VTL L=5e-08 W=5.4e-07 AD=7.56e-14 AS=6.3e-14 PD=1.36e-06 PS=1.36e-06 $X=2300 $Y=1960 $D=0
M20 20 A 19 VDD PMOS_VTL L=5e-08 W=5.4e-07 AD=7.695e-14 AS=7.56e-14 PD=1.365e-06 PS=1.36e-06 $X=2680 $Y=1960 $D=0
M21 13 CIN 20 VDD PMOS_VTL L=5e-08 W=5.4e-07 AD=6.3e-14 AS=7.695e-14 PD=1.36e-06 PS=1.365e-06 $X=3065 $Y=1960 $D=0
M22 14 11 13 VDD PMOS_VTL L=5e-08 W=3.6e-07 AD=5.13e-14 AS=6.3e-14 PD=1.005e-06 PS=1.36e-06 $X=3445 $Y=1960 $D=0
M23 VDD CIN 14 VDD PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=5.13e-14 PD=1e-06 PS=1.005e-06 $X=3830 $Y=1960 $D=0
M24 14 A VDD VDD PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=5.04e-14 PD=1e-06 PS=1e-06 $X=4210 $Y=1960 $D=0
M25 VDD B 14 VDD PMOS_VTL L=5e-08 W=3.6e-07 AD=4.14e-14 AS=5.04e-14 PD=9.5e-07 PS=1e-06 $X=4590 $Y=1960 $D=0
M26 COUT 11 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.07e-14 PD=5.9e-07 PS=5.9e-07 $X=5450 $Y=1960 $D=0
M27 SUM 13 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.07e-14 PD=5.9e-07 PS=5.9e-07 $X=6310 $Y=1960 $D=0
.ENDS
***************************************
.SUBCKT ICV_3 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
** N=26 EP=20 IP=36 FDC=112
X0 3 6 1 2 4 5 7 FullAdderMirror $T=0 0 0 0 $X=-50 $Y=-65
X1 10 6 8 9 11 5 12 FullAdderMirror $T=6800 6450 0 180 $X=-50 $Y=3170
X2 4 6 13 14 15 5 16 FullAdderMirror $T=6800 0 0 0 $X=6750 $Y=-65
X3 19 6 17 18 10 5 20 FullAdderMirror $T=13600 6450 0 180 $X=6750 $Y=3170
.ENDS
***************************************
.SUBCKT 16bitRCA GND SUM<15> SUM<7> A<8> VDD A<0> B<0> B<8> COUT CIN B<7> B<15> A<7> A<15> SUM<0> SUM<8> SUM<6> SUM<14> A<9> A<1>
+ B<1> B<9> B<6> B<14> A<6> A<14> SUM<1> SUM<9> SUM<5> SUM<13> A<10> A<2> B<10> B<2> B<13> B<5> A<5> A<13> SUM<2> SUM<10>
+ SUM<4> SUM<12> A<11> A<3> B<3> B<11> B<12> B<4> A<4> A<12> SUM<3> SUM<11>
** N=87 EP=52 IP=120 FDC=448
X4 A<0> B<0> CIN 2 GND VDD SUM<0> A<7> B<7> 4 1 SUM<7> A<1> B<1> 6 SUM<1> A<6> B<6> 8 SUM<6> ICV_3 $T=0 0 0 0 $X=-50 $Y=-65
X5 A<8> B<8> 1 3 GND VDD SUM<8> A<15> B<15> 5 COUT SUM<15> A<9> B<9> 7 SUM<9> A<14> B<14> 9 SUM<14> ICV_3 $T=0 6470 0 0 $X=-50 $Y=6405
X6 A<2> B<2> 6 10 GND VDD SUM<2> A<5> B<5> 12 8 SUM<5> A<3> B<3> 14 SUM<3> A<4> B<4> 14 SUM<4> ICV_3 $T=13600 0 0 0 $X=13550 $Y=-65
X7 A<10> B<10> 7 11 GND VDD SUM<10> A<13> B<13> 13 9 SUM<13> A<11> B<11> 15 SUM<11> A<12> B<12> 15 SUM<12> ICV_3 $T=13600 6470 0 0 $X=13550 $Y=6405
.ENDS
***************************************
