* SPICE NETLIST
***************************************

.SUBCKT M1_POLY_CDNS_586472688211
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT M2_M1_via
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_1
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_2
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT FullAdder Cin A B Cout GND VDD SUM
** N=25 EP=7 IP=31 FDC=28
M0 3 Cin GND GND NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.07e-14 PD=6.4e-07 PS=5.9e-07 $X=390 $Y=895 $D=1
M1 5 A 3 GND NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=770 $Y=895 $D=1
M2 3 B 5 GND NMOS_VTL L=5e-08 W=1.8e-07 AD=4.95e-14 AS=2.52e-14 PD=1.065e-06 PS=6.4e-07 $X=1150 $Y=895 $D=1
M3 23 A 3 GND NMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=4.95e-14 PD=1e-06 PS=1.065e-06 $X=1595 $Y=535 $D=1
M4 GND B 23 GND NMOS_VTL L=5e-08 W=3.6e-07 AD=4.14e-14 AS=5.04e-14 PD=9.5e-07 PS=1e-06 $X=1975 $Y=535 $D=1
M5 GND 5 7 GND NMOS_VTL L=5e-08 W=1.8e-07 AD=5.04e-14 AS=2.07e-14 PD=1.36e-06 PS=5.9e-07 $X=2855 $Y=895 $D=1
M6 24 A GND GND NMOS_VTL L=5e-08 W=5.4e-07 AD=7.56e-14 AS=5.04e-14 PD=1.36e-06 PS=1.36e-06 $X=3235 $Y=175 $D=1
M7 25 B 24 GND NMOS_VTL L=5e-08 W=5.4e-07 AD=7.56e-14 AS=7.56e-14 PD=1.36e-06 PS=1.36e-06 $X=3615 $Y=175 $D=1
M8 7 Cin 25 GND NMOS_VTL L=5e-08 W=5.4e-07 AD=5.04e-14 AS=7.56e-14 PD=1.36e-06 PS=1.36e-06 $X=3995 $Y=175 $D=1
M9 9 A 7 GND NMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=5.04e-14 PD=7.8e-07 PS=1.36e-06 $X=4375 $Y=895 $D=1
M10 7 B 9 GND NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=3.78e-14 PD=6.4e-07 PS=7.8e-07 $X=4895 $Y=895 $D=1
M11 9 Cin 7 GND NMOS_VTL L=5e-08 W=1.8e-07 AD=2.7e-14 AS=2.52e-14 PD=6.6e-07 PS=6.4e-07 $X=5275 $Y=895 $D=1
M12 Cout 5 GND GND NMOS_VTL L=5e-08 W=9e-08 AD=1.035e-14 AS=1.035e-14 PD=4.1e-07 PS=4.1e-07 $X=6225 $Y=1075 $D=1
M13 SUM 9 GND GND NMOS_VTL L=5e-08 W=9e-08 AD=1.035e-14 AS=1.035e-14 PD=4.1e-07 PS=4.1e-07 $X=7105 $Y=1075 $D=1
M14 VDD Cin 1 VDD PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=4.14e-14 PD=1e-06 PS=9.5e-07 $X=390 $Y=2675 $D=0
M15 20 A VDD VDD PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=5.04e-14 PD=1e-06 PS=1e-06 $X=770 $Y=2675 $D=0
M16 5 B 20 VDD PMOS_VTL L=5e-08 W=3.6e-07 AD=6.21e-14 AS=5.04e-14 PD=1.065e-06 PS=1e-06 $X=1150 $Y=2675 $D=0
M17 1 A 5 VDD PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=6.21e-14 PD=1e-06 PS=1.065e-06 $X=1595 $Y=2675 $D=0
M18 5 B 1 VDD PMOS_VTL L=5e-08 W=3.6e-07 AD=4.14e-14 AS=5.04e-14 PD=9.5e-07 PS=1e-06 $X=1975 $Y=2675 $D=0
M19 VDD 5 8 VDD PMOS_VTL L=5e-08 W=3.6e-07 AD=6.3e-14 AS=4.14e-14 PD=1.36e-06 PS=9.5e-07 $X=2855 $Y=2675 $D=0
M20 21 A VDD VDD PMOS_VTL L=5e-08 W=5.4e-07 AD=7.56e-14 AS=6.3e-14 PD=1.36e-06 PS=1.36e-06 $X=3235 $Y=2675 $D=0
M21 22 B 21 VDD PMOS_VTL L=5e-08 W=5.4e-07 AD=7.56e-14 AS=7.56e-14 PD=1.36e-06 PS=1.36e-06 $X=3615 $Y=2675 $D=0
M22 9 Cin 22 VDD PMOS_VTL L=5e-08 W=5.4e-07 AD=6.3e-14 AS=7.56e-14 PD=1.36e-06 PS=1.36e-06 $X=3995 $Y=2675 $D=0
M23 8 A 9 VDD PMOS_VTL L=5e-08 W=3.6e-07 AD=7.56e-14 AS=6.3e-14 PD=1.14e-06 PS=1.36e-06 $X=4375 $Y=2675 $D=0
M24 9 B 8 VDD PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=7.56e-14 PD=1e-06 PS=1.14e-06 $X=4895 $Y=2675 $D=0
M25 8 Cin 9 VDD PMOS_VTL L=5e-08 W=3.6e-07 AD=5.4e-14 AS=5.04e-14 PD=1.02e-06 PS=1e-06 $X=5275 $Y=2675 $D=0
M26 Cout 5 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.07e-14 PD=5.9e-07 PS=5.9e-07 $X=6225 $Y=2675 $D=0
M27 SUM 9 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.07e-14 PD=5.9e-07 PS=5.9e-07 $X=7105 $Y=2675 $D=0
.ENDS
***************************************
