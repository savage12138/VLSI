* SPICE NETLIST
***************************************

.SUBCKT M1_POLY_CDNS_586656140050
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT M2_M1_via
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT FullAdderMirror CIN A B COUT GND VDD SUM
** N=24 EP=7 IP=19 FDC=28
M0 GND A 1 GND NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.07e-14 PD=6.4e-07 PS=5.9e-07 $X=890 $Y=355 $D=1
M1 22 A GND GND NMOS_VTL L=5e-08 W=1.8e-07 AD=2.565e-14 AS=2.52e-14 PD=6.45e-07 PS=6.4e-07 $X=1270 $Y=355 $D=1
M2 3 B 22 GND NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.565e-14 PD=6.4e-07 PS=6.45e-07 $X=1655 $Y=355 $D=1
M3 1 CIN 3 GND NMOS_VTL L=5e-08 W=1.8e-07 AD=2.565e-14 AS=2.52e-14 PD=6.45e-07 PS=6.4e-07 $X=2035 $Y=355 $D=1
M4 GND B 1 GND NMOS_VTL L=5e-08 W=1.8e-07 AD=3.15e-14 AS=2.565e-14 PD=8.2e-07 PS=6.45e-07 $X=2420 $Y=355 $D=1
M5 23 B GND GND NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=3.15e-14 PD=8.2e-07 PS=8.2e-07 $X=2800 $Y=175 $D=1
M6 24 A 23 GND NMOS_VTL L=5e-08 W=2.7e-07 AD=3.8475e-14 AS=3.78e-14 PD=8.25e-07 PS=8.2e-07 $X=3180 $Y=175 $D=1
M7 7 CIN 24 GND NMOS_VTL L=5e-08 W=2.7e-07 AD=3.15e-14 AS=3.8475e-14 PD=8.2e-07 PS=8.25e-07 $X=3565 $Y=175 $D=1
M8 8 3 7 GND NMOS_VTL L=5e-08 W=1.8e-07 AD=2.565e-14 AS=3.15e-14 PD=6.45e-07 PS=8.2e-07 $X=3945 $Y=355 $D=1
M9 GND CIN 8 GND NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.565e-14 PD=6.4e-07 PS=6.45e-07 $X=4330 $Y=355 $D=1
M10 8 A GND GND NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=4710 $Y=355 $D=1
M11 GND B 8 GND NMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.52e-14 PD=5.9e-07 PS=6.4e-07 $X=5090 $Y=355 $D=1
M12 COUT 3 GND GND NMOS_VTL L=5e-08 W=9e-08 AD=1.035e-14 AS=1.035e-14 PD=4.1e-07 PS=4.1e-07 $X=5950 $Y=535 $D=1
M13 SUM 7 GND GND NMOS_VTL L=5e-08 W=9e-08 AD=1.035e-14 AS=1.035e-14 PD=4.1e-07 PS=4.1e-07 $X=6810 $Y=535 $D=1
M14 VDD A 4 VDD PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=4.14e-14 PD=1e-06 PS=9.5e-07 $X=890 $Y=1960 $D=0
M15 19 A VDD VDD PMOS_VTL L=5e-08 W=3.6e-07 AD=5.13e-14 AS=5.04e-14 PD=1.005e-06 PS=1e-06 $X=1270 $Y=1960 $D=0
M16 3 B 19 VDD PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=5.13e-14 PD=1e-06 PS=1.005e-06 $X=1655 $Y=1960 $D=0
M17 4 CIN 3 VDD PMOS_VTL L=5e-08 W=3.6e-07 AD=5.13e-14 AS=5.04e-14 PD=1.005e-06 PS=1e-06 $X=2035 $Y=1960 $D=0
M18 VDD B 4 VDD PMOS_VTL L=5e-08 W=3.6e-07 AD=6.3e-14 AS=5.13e-14 PD=1.36e-06 PS=1.005e-06 $X=2420 $Y=1960 $D=0
M19 20 B VDD VDD PMOS_VTL L=5e-08 W=5.4e-07 AD=7.56e-14 AS=6.3e-14 PD=1.36e-06 PS=1.36e-06 $X=2800 $Y=1960 $D=0
M20 21 A 20 VDD PMOS_VTL L=5e-08 W=5.4e-07 AD=7.695e-14 AS=7.56e-14 PD=1.365e-06 PS=1.36e-06 $X=3180 $Y=1960 $D=0
M21 7 CIN 21 VDD PMOS_VTL L=5e-08 W=5.4e-07 AD=6.3e-14 AS=7.695e-14 PD=1.36e-06 PS=1.365e-06 $X=3565 $Y=1960 $D=0
M22 9 3 7 VDD PMOS_VTL L=5e-08 W=3.6e-07 AD=5.13e-14 AS=6.3e-14 PD=1.005e-06 PS=1.36e-06 $X=3945 $Y=1960 $D=0
M23 VDD CIN 9 VDD PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=5.13e-14 PD=1e-06 PS=1.005e-06 $X=4330 $Y=1960 $D=0
M24 9 A VDD VDD PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=5.04e-14 PD=1e-06 PS=1e-06 $X=4710 $Y=1960 $D=0
M25 VDD B 9 VDD PMOS_VTL L=5e-08 W=3.6e-07 AD=4.14e-14 AS=5.04e-14 PD=9.5e-07 PS=1e-06 $X=5090 $Y=1960 $D=0
M26 COUT 3 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.07e-14 PD=5.9e-07 PS=5.9e-07 $X=5950 $Y=1960 $D=0
M27 SUM 7 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.07e-14 PD=5.9e-07 PS=5.9e-07 $X=6810 $Y=1960 $D=0
.ENDS
***************************************
